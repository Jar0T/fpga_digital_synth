--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.common_pkg.all;

package osc_pkg is

    constant PHASE_WIDTH : integer := 32;
    constant SAMPLE_WIDTH : integer := 16;
    constant SAMPLE_ADDR_WIDTH : integer := 9;
    
    type t_phase_step_array is array(0 to N_CHANNELS - 1) of unsigned(PHASE_WIDTH - 1 downto 0);
    type t_sample_array is array(0 to N_CHANNELS - 1) of signed(SAMPLE_WIDTH - 1 downto 0);
    
    type t_wave_lut is array(0 to 2**SAMPLE_ADDR_WIDTH - 1) of signed(SAMPLE_WIDTH - 1 downto 0);
    
    constant SINE_WAVE_INIT : t_wave_lut;

end osc_pkg;

package body osc_pkg is

    constant SINE_WAVE_INIT : t_wave_lut := (
        0 => to_signed(0, 16),
        1 => to_signed(402, 16),
        2 => to_signed(804, 16),
        3 => to_signed(1206, 16),
        4 => to_signed(1607, 16),
        5 => to_signed(2009, 16),
        6 => to_signed(2410, 16),
        7 => to_signed(2811, 16),
        8 => to_signed(3211, 16),
        9 => to_signed(3611, 16),
        10 => to_signed(4011, 16),
        11 => to_signed(4409, 16),
        12 => to_signed(4807, 16),
        13 => to_signed(5205, 16),
        14 => to_signed(5601, 16),
        15 => to_signed(5997, 16),
        16 => to_signed(6392, 16),
        17 => to_signed(6786, 16),
        18 => to_signed(7179, 16),
        19 => to_signed(7571, 16),
        20 => to_signed(7961, 16),
        21 => to_signed(8351, 16),
        22 => to_signed(8739, 16),
        23 => to_signed(9126, 16),
        24 => to_signed(9511, 16),
        25 => to_signed(9895, 16),
        26 => to_signed(10278, 16),
        27 => to_signed(10659, 16),
        28 => to_signed(11038, 16),
        29 => to_signed(11416, 16),
        30 => to_signed(11792, 16),
        31 => to_signed(12166, 16),
        32 => to_signed(12539, 16),
        33 => to_signed(12909, 16),
        34 => to_signed(13278, 16),
        35 => to_signed(13645, 16),
        36 => to_signed(14009, 16),
        37 => to_signed(14372, 16),
        38 => to_signed(14732, 16),
        39 => to_signed(15090, 16),
        40 => to_signed(15446, 16),
        41 => to_signed(15799, 16),
        42 => to_signed(16150, 16),
        43 => to_signed(16499, 16),
        44 => to_signed(16845, 16),
        45 => to_signed(17189, 16),
        46 => to_signed(17530, 16),
        47 => to_signed(17868, 16),
        48 => to_signed(18204, 16),
        49 => to_signed(18537, 16),
        50 => to_signed(18867, 16),
        51 => to_signed(19194, 16),
        52 => to_signed(19519, 16),
        53 => to_signed(19840, 16),
        54 => to_signed(20159, 16),
        55 => to_signed(20474, 16),
        56 => to_signed(20787, 16),
        57 => to_signed(21096, 16),
        58 => to_signed(21402, 16),
        59 => to_signed(21705, 16),
        60 => to_signed(22004, 16),
        61 => to_signed(22301, 16),
        62 => to_signed(22594, 16),
        63 => to_signed(22883, 16),
        64 => to_signed(23169, 16),
        65 => to_signed(23452, 16),
        66 => to_signed(23731, 16),
        67 => to_signed(24006, 16),
        68 => to_signed(24278, 16),
        69 => to_signed(24546, 16),
        70 => to_signed(24811, 16),
        71 => to_signed(25072, 16),
        72 => to_signed(25329, 16),
        73 => to_signed(25582, 16),
        74 => to_signed(25831, 16),
        75 => to_signed(26077, 16),
        76 => to_signed(26318, 16),
        77 => to_signed(26556, 16),
        78 => to_signed(26789, 16),
        79 => to_signed(27019, 16),
        80 => to_signed(27244, 16),
        81 => to_signed(27466, 16),
        82 => to_signed(27683, 16),
        83 => to_signed(27896, 16),
        84 => to_signed(28105, 16),
        85 => to_signed(28309, 16),
        86 => to_signed(28510, 16),
        87 => to_signed(28706, 16),
        88 => to_signed(28897, 16),
        89 => to_signed(29085, 16),
        90 => to_signed(29268, 16),
        91 => to_signed(29446, 16),
        92 => to_signed(29621, 16),
        93 => to_signed(29790, 16),
        94 => to_signed(29955, 16),
        95 => to_signed(30116, 16),
        96 => to_signed(30272, 16),
        97 => to_signed(30424, 16),
        98 => to_signed(30571, 16),
        99 => to_signed(30713, 16),
        100 => to_signed(30851, 16),
        101 => to_signed(30984, 16),
        102 => to_signed(31113, 16),
        103 => to_signed(31236, 16),
        104 => to_signed(31356, 16),
        105 => to_signed(31470, 16),
        106 => to_signed(31580, 16),
        107 => to_signed(31684, 16),
        108 => to_signed(31785, 16),
        109 => to_signed(31880, 16),
        110 => to_signed(31970, 16),
        111 => to_signed(32056, 16),
        112 => to_signed(32137, 16),
        113 => to_signed(32213, 16),
        114 => to_signed(32284, 16),
        115 => to_signed(32350, 16),
        116 => to_signed(32412, 16),
        117 => to_signed(32468, 16),
        118 => to_signed(32520, 16),
        119 => to_signed(32567, 16),
        120 => to_signed(32609, 16),
        121 => to_signed(32646, 16),
        122 => to_signed(32678, 16),
        123 => to_signed(32705, 16),
        124 => to_signed(32727, 16),
        125 => to_signed(32744, 16),
        126 => to_signed(32757, 16),
        127 => to_signed(32764, 16),
        128 => to_signed(32767, 16),
        129 => to_signed(32764, 16),
        130 => to_signed(32757, 16),
        131 => to_signed(32744, 16),
        132 => to_signed(32727, 16),
        133 => to_signed(32705, 16),
        134 => to_signed(32678, 16),
        135 => to_signed(32646, 16),
        136 => to_signed(32609, 16),
        137 => to_signed(32567, 16),
        138 => to_signed(32520, 16),
        139 => to_signed(32468, 16),
        140 => to_signed(32412, 16),
        141 => to_signed(32350, 16),
        142 => to_signed(32284, 16),
        143 => to_signed(32213, 16),
        144 => to_signed(32137, 16),
        145 => to_signed(32056, 16),
        146 => to_signed(31970, 16),
        147 => to_signed(31880, 16),
        148 => to_signed(31785, 16),
        149 => to_signed(31684, 16),
        150 => to_signed(31580, 16),
        151 => to_signed(31470, 16),
        152 => to_signed(31356, 16),
        153 => to_signed(31236, 16),
        154 => to_signed(31113, 16),
        155 => to_signed(30984, 16),
        156 => to_signed(30851, 16),
        157 => to_signed(30713, 16),
        158 => to_signed(30571, 16),
        159 => to_signed(30424, 16),
        160 => to_signed(30272, 16),
        161 => to_signed(30116, 16),
        162 => to_signed(29955, 16),
        163 => to_signed(29790, 16),
        164 => to_signed(29621, 16),
        165 => to_signed(29446, 16),
        166 => to_signed(29268, 16),
        167 => to_signed(29085, 16),
        168 => to_signed(28897, 16),
        169 => to_signed(28706, 16),
        170 => to_signed(28510, 16),
        171 => to_signed(28309, 16),
        172 => to_signed(28105, 16),
        173 => to_signed(27896, 16),
        174 => to_signed(27683, 16),
        175 => to_signed(27466, 16),
        176 => to_signed(27244, 16),
        177 => to_signed(27019, 16),
        178 => to_signed(26789, 16),
        179 => to_signed(26556, 16),
        180 => to_signed(26318, 16),
        181 => to_signed(26077, 16),
        182 => to_signed(25831, 16),
        183 => to_signed(25582, 16),
        184 => to_signed(25329, 16),
        185 => to_signed(25072, 16),
        186 => to_signed(24811, 16),
        187 => to_signed(24546, 16),
        188 => to_signed(24278, 16),
        189 => to_signed(24006, 16),
        190 => to_signed(23731, 16),
        191 => to_signed(23452, 16),
        192 => to_signed(23169, 16),
        193 => to_signed(22883, 16),
        194 => to_signed(22594, 16),
        195 => to_signed(22301, 16),
        196 => to_signed(22004, 16),
        197 => to_signed(21705, 16),
        198 => to_signed(21402, 16),
        199 => to_signed(21096, 16),
        200 => to_signed(20787, 16),
        201 => to_signed(20474, 16),
        202 => to_signed(20159, 16),
        203 => to_signed(19840, 16),
        204 => to_signed(19519, 16),
        205 => to_signed(19194, 16),
        206 => to_signed(18867, 16),
        207 => to_signed(18537, 16),
        208 => to_signed(18204, 16),
        209 => to_signed(17868, 16),
        210 => to_signed(17530, 16),
        211 => to_signed(17189, 16),
        212 => to_signed(16845, 16),
        213 => to_signed(16499, 16),
        214 => to_signed(16150, 16),
        215 => to_signed(15799, 16),
        216 => to_signed(15446, 16),
        217 => to_signed(15090, 16),
        218 => to_signed(14732, 16),
        219 => to_signed(14372, 16),
        220 => to_signed(14009, 16),
        221 => to_signed(13645, 16),
        222 => to_signed(13278, 16),
        223 => to_signed(12909, 16),
        224 => to_signed(12539, 16),
        225 => to_signed(12166, 16),
        226 => to_signed(11792, 16),
        227 => to_signed(11416, 16),
        228 => to_signed(11038, 16),
        229 => to_signed(10659, 16),
        230 => to_signed(10278, 16),
        231 => to_signed(9895, 16),
        232 => to_signed(9511, 16),
        233 => to_signed(9126, 16),
        234 => to_signed(8739, 16),
        235 => to_signed(8351, 16),
        236 => to_signed(7961, 16),
        237 => to_signed(7571, 16),
        238 => to_signed(7179, 16),
        239 => to_signed(6786, 16),
        240 => to_signed(6392, 16),
        241 => to_signed(5997, 16),
        242 => to_signed(5601, 16),
        243 => to_signed(5205, 16),
        244 => to_signed(4807, 16),
        245 => to_signed(4409, 16),
        246 => to_signed(4011, 16),
        247 => to_signed(3611, 16),
        248 => to_signed(3211, 16),
        249 => to_signed(2811, 16),
        250 => to_signed(2410, 16),
        251 => to_signed(2009, 16),
        252 => to_signed(1607, 16),
        253 => to_signed(1206, 16),
        254 => to_signed(804, 16),
        255 => to_signed(402, 16),
        256 => to_signed(0, 16),
        257 => to_signed(-402, 16),
        258 => to_signed(-804, 16),
        259 => to_signed(-1206, 16),
        260 => to_signed(-1607, 16),
        261 => to_signed(-2009, 16),
        262 => to_signed(-2410, 16),
        263 => to_signed(-2811, 16),
        264 => to_signed(-3211, 16),
        265 => to_signed(-3611, 16),
        266 => to_signed(-4011, 16),
        267 => to_signed(-4409, 16),
        268 => to_signed(-4807, 16),
        269 => to_signed(-5205, 16),
        270 => to_signed(-5601, 16),
        271 => to_signed(-5997, 16),
        272 => to_signed(-6392, 16),
        273 => to_signed(-6786, 16),
        274 => to_signed(-7179, 16),
        275 => to_signed(-7571, 16),
        276 => to_signed(-7961, 16),
        277 => to_signed(-8351, 16),
        278 => to_signed(-8739, 16),
        279 => to_signed(-9126, 16),
        280 => to_signed(-9511, 16),
        281 => to_signed(-9895, 16),
        282 => to_signed(-10278, 16),
        283 => to_signed(-10659, 16),
        284 => to_signed(-11038, 16),
        285 => to_signed(-11416, 16),
        286 => to_signed(-11792, 16),
        287 => to_signed(-12166, 16),
        288 => to_signed(-12539, 16),
        289 => to_signed(-12909, 16),
        290 => to_signed(-13278, 16),
        291 => to_signed(-13645, 16),
        292 => to_signed(-14009, 16),
        293 => to_signed(-14372, 16),
        294 => to_signed(-14732, 16),
        295 => to_signed(-15090, 16),
        296 => to_signed(-15446, 16),
        297 => to_signed(-15799, 16),
        298 => to_signed(-16150, 16),
        299 => to_signed(-16499, 16),
        300 => to_signed(-16845, 16),
        301 => to_signed(-17189, 16),
        302 => to_signed(-17530, 16),
        303 => to_signed(-17868, 16),
        304 => to_signed(-18204, 16),
        305 => to_signed(-18537, 16),
        306 => to_signed(-18867, 16),
        307 => to_signed(-19194, 16),
        308 => to_signed(-19519, 16),
        309 => to_signed(-19840, 16),
        310 => to_signed(-20159, 16),
        311 => to_signed(-20474, 16),
        312 => to_signed(-20787, 16),
        313 => to_signed(-21096, 16),
        314 => to_signed(-21402, 16),
        315 => to_signed(-21705, 16),
        316 => to_signed(-22004, 16),
        317 => to_signed(-22301, 16),
        318 => to_signed(-22594, 16),
        319 => to_signed(-22883, 16),
        320 => to_signed(-23169, 16),
        321 => to_signed(-23452, 16),
        322 => to_signed(-23731, 16),
        323 => to_signed(-24006, 16),
        324 => to_signed(-24278, 16),
        325 => to_signed(-24546, 16),
        326 => to_signed(-24811, 16),
        327 => to_signed(-25072, 16),
        328 => to_signed(-25329, 16),
        329 => to_signed(-25582, 16),
        330 => to_signed(-25831, 16),
        331 => to_signed(-26077, 16),
        332 => to_signed(-26318, 16),
        333 => to_signed(-26556, 16),
        334 => to_signed(-26789, 16),
        335 => to_signed(-27019, 16),
        336 => to_signed(-27244, 16),
        337 => to_signed(-27466, 16),
        338 => to_signed(-27683, 16),
        339 => to_signed(-27896, 16),
        340 => to_signed(-28105, 16),
        341 => to_signed(-28309, 16),
        342 => to_signed(-28510, 16),
        343 => to_signed(-28706, 16),
        344 => to_signed(-28897, 16),
        345 => to_signed(-29085, 16),
        346 => to_signed(-29268, 16),
        347 => to_signed(-29446, 16),
        348 => to_signed(-29621, 16),
        349 => to_signed(-29790, 16),
        350 => to_signed(-29955, 16),
        351 => to_signed(-30116, 16),
        352 => to_signed(-30272, 16),
        353 => to_signed(-30424, 16),
        354 => to_signed(-30571, 16),
        355 => to_signed(-30713, 16),
        356 => to_signed(-30851, 16),
        357 => to_signed(-30984, 16),
        358 => to_signed(-31113, 16),
        359 => to_signed(-31236, 16),
        360 => to_signed(-31356, 16),
        361 => to_signed(-31470, 16),
        362 => to_signed(-31580, 16),
        363 => to_signed(-31684, 16),
        364 => to_signed(-31785, 16),
        365 => to_signed(-31880, 16),
        366 => to_signed(-31970, 16),
        367 => to_signed(-32056, 16),
        368 => to_signed(-32137, 16),
        369 => to_signed(-32213, 16),
        370 => to_signed(-32284, 16),
        371 => to_signed(-32350, 16),
        372 => to_signed(-32412, 16),
        373 => to_signed(-32468, 16),
        374 => to_signed(-32520, 16),
        375 => to_signed(-32567, 16),
        376 => to_signed(-32609, 16),
        377 => to_signed(-32646, 16),
        378 => to_signed(-32678, 16),
        379 => to_signed(-32705, 16),
        380 => to_signed(-32727, 16),
        381 => to_signed(-32744, 16),
        382 => to_signed(-32757, 16),
        383 => to_signed(-32764, 16),
        384 => to_signed(-32767, 16),
        385 => to_signed(-32764, 16),
        386 => to_signed(-32757, 16),
        387 => to_signed(-32744, 16),
        388 => to_signed(-32727, 16),
        389 => to_signed(-32705, 16),
        390 => to_signed(-32678, 16),
        391 => to_signed(-32646, 16),
        392 => to_signed(-32609, 16),
        393 => to_signed(-32567, 16),
        394 => to_signed(-32520, 16),
        395 => to_signed(-32468, 16),
        396 => to_signed(-32412, 16),
        397 => to_signed(-32350, 16),
        398 => to_signed(-32284, 16),
        399 => to_signed(-32213, 16),
        400 => to_signed(-32137, 16),
        401 => to_signed(-32056, 16),
        402 => to_signed(-31970, 16),
        403 => to_signed(-31880, 16),
        404 => to_signed(-31785, 16),
        405 => to_signed(-31684, 16),
        406 => to_signed(-31580, 16),
        407 => to_signed(-31470, 16),
        408 => to_signed(-31356, 16),
        409 => to_signed(-31236, 16),
        410 => to_signed(-31113, 16),
        411 => to_signed(-30984, 16),
        412 => to_signed(-30851, 16),
        413 => to_signed(-30713, 16),
        414 => to_signed(-30571, 16),
        415 => to_signed(-30424, 16),
        416 => to_signed(-30272, 16),
        417 => to_signed(-30116, 16),
        418 => to_signed(-29955, 16),
        419 => to_signed(-29790, 16),
        420 => to_signed(-29621, 16),
        421 => to_signed(-29446, 16),
        422 => to_signed(-29268, 16),
        423 => to_signed(-29085, 16),
        424 => to_signed(-28897, 16),
        425 => to_signed(-28706, 16),
        426 => to_signed(-28510, 16),
        427 => to_signed(-28309, 16),
        428 => to_signed(-28105, 16),
        429 => to_signed(-27896, 16),
        430 => to_signed(-27683, 16),
        431 => to_signed(-27466, 16),
        432 => to_signed(-27244, 16),
        433 => to_signed(-27019, 16),
        434 => to_signed(-26789, 16),
        435 => to_signed(-26556, 16),
        436 => to_signed(-26318, 16),
        437 => to_signed(-26077, 16),
        438 => to_signed(-25831, 16),
        439 => to_signed(-25582, 16),
        440 => to_signed(-25329, 16),
        441 => to_signed(-25072, 16),
        442 => to_signed(-24811, 16),
        443 => to_signed(-24546, 16),
        444 => to_signed(-24278, 16),
        445 => to_signed(-24006, 16),
        446 => to_signed(-23731, 16),
        447 => to_signed(-23452, 16),
        448 => to_signed(-23169, 16),
        449 => to_signed(-22883, 16),
        450 => to_signed(-22594, 16),
        451 => to_signed(-22301, 16),
        452 => to_signed(-22004, 16),
        453 => to_signed(-21705, 16),
        454 => to_signed(-21402, 16),
        455 => to_signed(-21096, 16),
        456 => to_signed(-20787, 16),
        457 => to_signed(-20474, 16),
        458 => to_signed(-20159, 16),
        459 => to_signed(-19840, 16),
        460 => to_signed(-19519, 16),
        461 => to_signed(-19194, 16),
        462 => to_signed(-18867, 16),
        463 => to_signed(-18537, 16),
        464 => to_signed(-18204, 16),
        465 => to_signed(-17868, 16),
        466 => to_signed(-17530, 16),
        467 => to_signed(-17189, 16),
        468 => to_signed(-16845, 16),
        469 => to_signed(-16499, 16),
        470 => to_signed(-16150, 16),
        471 => to_signed(-15799, 16),
        472 => to_signed(-15446, 16),
        473 => to_signed(-15090, 16),
        474 => to_signed(-14732, 16),
        475 => to_signed(-14372, 16),
        476 => to_signed(-14009, 16),
        477 => to_signed(-13645, 16),
        478 => to_signed(-13278, 16),
        479 => to_signed(-12909, 16),
        480 => to_signed(-12539, 16),
        481 => to_signed(-12166, 16),
        482 => to_signed(-11792, 16),
        483 => to_signed(-11416, 16),
        484 => to_signed(-11038, 16),
        485 => to_signed(-10659, 16),
        486 => to_signed(-10278, 16),
        487 => to_signed(-9895, 16),
        488 => to_signed(-9511, 16),
        489 => to_signed(-9126, 16),
        490 => to_signed(-8739, 16),
        491 => to_signed(-8351, 16),
        492 => to_signed(-7961, 16),
        493 => to_signed(-7571, 16),
        494 => to_signed(-7179, 16),
        495 => to_signed(-6786, 16),
        496 => to_signed(-6392, 16),
        497 => to_signed(-5997, 16),
        498 => to_signed(-5601, 16),
        499 => to_signed(-5205, 16),
        500 => to_signed(-4807, 16),
        501 => to_signed(-4409, 16),
        502 => to_signed(-4011, 16),
        503 => to_signed(-3611, 16),
        504 => to_signed(-3211, 16),
        505 => to_signed(-2811, 16),
        506 => to_signed(-2410, 16),
        507 => to_signed(-2009, 16),
        508 => to_signed(-1607, 16),
        509 => to_signed(-1206, 16),
        510 => to_signed(-804, 16),
        511 => to_signed(-402, 16)
    );
 
end osc_pkg;
